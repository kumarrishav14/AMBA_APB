`include "uvm_macros.svh"
`include "interface.sv"
`include "config_objs.svh"
`include "transaction.sv"
`include "rnd_sequence.sv"
`include "driver.sv"
`include "monitor.sv"
`include "fun_cov.sv"
`include "agent.sv"
`include "test.sv"