`include "uvm_macros.svh"
`include "interface.sv"
`include "transaction.sv"
`include "rnd_sequence.sv"
`include "driver.sv"
`include "monitor.sv"
`include "agent.sv"