`include "generator.sv"
`include "driver.sv"
`include "ip_monitor.sv"
`include "op_monitor.sv"
`include "ref_model.sv"
`include "scoreboard.sv"
`include "environment.sv"
`include "test.sv"
`include "interface.sv"
