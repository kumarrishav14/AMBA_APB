class ref_model;
    mailbox #(transaction) ipmon2rm;
    mailbox #(transaction) rm2sb;

    const int ram_depth = 2**4;
    // Memory for 4KB RAM
    bit [31:0] ram_mem [];

    transaction trans, trans2sb;
    function new(mailbox #(transaction) ipmon2rm, mailbox #(transaction) rm2sb);
        this.ipmon2rm = ipmon2rm;
        this.rm2sb = rm2sb;

        trans = new;
        ram_mem = new[ram_depth];
    endfunction //new()

    
    
    task gen_op();
        for(int i=0; i<trans.PADDR.size(); i++) begin
            if(trans.PRESETn == 0) begin
                continue;
            end
            if(trans.PADDR[i] >= ram_depth) begin
                trans.PSLVERR = 1;
                trans.PRDATA[i] = 32'b0;
                trans.PREADY = 1;
                continue;
            end

            if(trans.PWRITE == 1) begin
                ram_mem [trans.PADDR[i]] = trans.PWDATA[i];
                trans.PRDATA[i] = 32'b0;
                trans.PREADY = 1;
                trans.PSLVERR = 0;
            end
            else begin
                trans.PRDATA[i] = ram_mem [trans.PADDR[i]];
                trans.PREADY = 1;
                trans.PSLVERR = 0;
            end
                

        end
    endtask //gen_op

    task start();
        fork
            forever begin
                ipmon2rm.get(trans);
                gen_op();
                trans2sb = new trans;
                //trans2sb.printf("OUTPUT GENERATED BY RM");
                rm2sb.put(trans2sb);
            end
        join_none
    endtask //start
endclass //ref_model